*MOSIS 2U CMOS MODELS

.MODEL nfet NMOS LEVEL=2 LD=0.115U TOX=423E-10
+NSUB=1.0125225E+16 VTO=0.822163 KP=4.893760E-5 GAMMA=0.47
+PHI=0.6 UO=599.496 UEXP=5.324966E-3 UCRIT=12714.2
+DELTA=3.39718E-5 VMAX=65466.1 XJ=0.55U LAMBDA=1.991479e-2
+NFS=5.666758E+11 NEFF=1.0010E-2 NSS=0.0 TPG=1.00
+RSH=0 CGSO=0.9388E-10 CGDO=0.9388E-10 CJ=1.4563E-4
+MJ=0.6 CJSW=6.617E-10 MJSW=0.31

.MODEL pfet PMOS LEVEL=2 LD=0.18U TOX=423E-10
+NSUB=1.421645E+15 VTO=-0.776658 KP=1.916950E-5 GAMMA=0.52
+PHI=0.6 UO=234.831 UEXP=0.142293 UCRIT=20967
+DELTA=1.0E-6 VMAX=34600.2 XJ=0.41U LAMBDA=4.921086E-2
+NFS=4.744781E+11 NEFF=1.0010E-2 NSS=0.0 TPG=-1.00
+RSH=0 CGSO=1.469E-10 CGDO=1.469E-10 CJ=2.4E-4
+MJ=0.5 CJSW=3.62E-10 MJSW=0.29
